`ifndef UARTSTATES
`define UARTSTATES
/*
 Universidade Estadual de Feira de Santana
 TEC499 - MI - Sistemas Digitais

 States used on UART's Rx and Tx modules

*/

/*ALU Operations*/
`define IDLE  2'b00
`define START 2'b01
`define WORK 2'b10
`define STOP 2'b11

`endif //UARTSTATES
